`default_nettype none

module Main;
   initial begin 
      $display("Hello, World!"); 
      $finish;
   end
endmodule
